module algo (clock, in1, in2, in3, past_data, out);
   input wire in1, in2, in3;
   input wire [31:0] past_data;
   output reg out;

   reg result;

   always @(posedge clock) begin
      // use a complex algorithm to set reg result based on in1, in2, in3, and past_data
      out = result;
   end
endmodule